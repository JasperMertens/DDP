`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    10:29:29 11/14/2016 
// Design Name: 
// Module Name:    compute_ddp_wrapper 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module compute_ddp_wrapper(clk, rst, a0, a1, b0, b1, result, result_ready);
input clk;
input rst;
input [3:0] a0, a1, b0, b1;

output [4:0] result;		// in this example, result is a0+b0 and then a1+b1 
output result_ready;		// goes high when a0+b0 is computed and a1+b1 is computed

wire [3:0] ma_out, mb_out;
wire [4:0] compute_out;


// control signals generated by the FSM
reg ma_sel, mb_sel, compute_start, result_ready;

// control signals read by the FSM
wire compute_done;

// state variables
reg [2:0] state, nextstate;


//// ALU is described here

// Description of compute_ddp is in the other file.
// Description of mux2x1 is at the bottom of this file.
mux2x1 ma(.in0(a0), .in1(a1), .sel(ma_sel), .out(ma_out));
mux2x1 mb(.in0(b0), .in1(b1), .sel(mb_sel), .out(mb_out));
compute_ddp	compute( .clk(clk), .rst(rst), .start(compute_start), .a(ma_out), .b(mb_out), .c(compute_out), .done(compute_done) );
assign result = compute_out;

//// FSM is described here

always @(posedge clk)
begin
	if(rst)	// outside reset brings the FSM to init state (i.e. state0)
 		state <= 3'd0;
	else
		state <= nextstate;
end		

always @(*)
begin
	case(state)
	3'd0: begin		// Initial idle state
				ma_sel<=1'b0; mb_sel<=1'b0; compute_start<=1'b0; result_ready<=1'b0;
			end

	3'd1: begin		// initiate computation of a0+b0
				ma_sel<=1'b0; mb_sel<=1'b0; compute_start<=1'b1; result_ready<=1'b0;
			end
	3'd2: begin		// wait for this computation to finish
				ma_sel<=1'b0; mb_sel<=1'b0; compute_start<=1'b0; result_ready<=1'b0;
			end
	3'd3: begin		// set result_ready
				ma_sel<=1'b0; mb_sel<=1'b0; compute_start<=1'b0; result_ready<=1'b1;
			end

			
	3'd4: begin		// then initiate computation of a1+b1
				ma_sel<=1'b1; mb_sel<=1'b1; compute_start<=1'b1; result_ready<=1'b0;
			end
	3'd5: begin		// again wait for this computation to finish
				ma_sel<=1'b1; mb_sel<=1'b1; compute_start<=1'b0; result_ready<=1'b0;
			end			
	3'd6: begin		// set result_ready
				ma_sel<=1'b1; mb_sel<=1'b1; compute_start<=1'b0; result_ready<=1'b1;
			end			

	3'd7: begin		// END: no work 
				ma_sel<=1'b0; mb_sel<=1'b0; compute_start<=1'b0; result_ready<=1'b0;
			end
	default: begin		
				ma_sel<=1'b0; mb_sel<=1'b0; compute_start<=1'b0; result_ready<=1'b0;
			end
	endcase
end


// nextstate logic
always @(*)
begin
	case(state)
	3'd0: nextstate <=3'd1;

	3'd1: nextstate <=3'd2;		// initiates a0+b0
	3'd2: begin
				if(compute_done)	// wait for the computation to finish
					nextstate <=3'd3;
				else
					nextstate <=3'd2;
			end		
	3'd3: nextstate <=3'd4;		

	3'd4: nextstate <=3'd5;		// initiates a1+b1
	3'd5: begin
				if(compute_done)	// wait for the computation to finish
					nextstate <=3'd6;
				else
					nextstate <=3'd5;
			end		
	3'd6: nextstate <=3'd7;

	3'd7: nextstate <=3'd7;		// FSM halts here
	default: nextstate <=3'd0;	
	endcase
end	
	
endmodule



module mux2x1(in0, in1, sel, out);
input [3:0] in0, in1;
input sel;
output [3:0] out;

assign out = (sel==1'b0) ? in0 : in1;

endmodule

